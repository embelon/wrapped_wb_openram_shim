VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_wb_openram_shim
  CLASS BLOCK ;
  FOREIGN wrapped_wb_openram_shim ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 28.600 40.000 29.200 ;
    END
  END active
  PIN openram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 296.520 40.000 297.120 ;
    END
  END openram_addr0[0]
  PIN openram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END openram_addr0[1]
  PIN openram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END openram_addr0[2]
  PIN openram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END openram_addr0[3]
  PIN openram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 93.880 40.000 94.480 ;
    END
  END openram_addr0[4]
  PIN openram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END openram_addr0[5]
  PIN openram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END openram_addr0[6]
  PIN openram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 141.480 40.000 142.080 ;
    END
  END openram_addr0[7]
  PIN openram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END openram_clk0
  PIN openram_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 164.600 40.000 165.200 ;
    END
  END openram_csb0
  PIN openram_din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 102.040 40.000 102.640 ;
    END
  END openram_din0[0]
  PIN openram_din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END openram_din0[10]
  PIN openram_din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END openram_din0[11]
  PIN openram_din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END openram_din0[12]
  PIN openram_din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END openram_din0[13]
  PIN openram_din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END openram_din0[14]
  PIN openram_din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END openram_din0[15]
  PIN openram_din0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END openram_din0[16]
  PIN openram_din0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END openram_din0[17]
  PIN openram_din0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 59.880 40.000 60.480 ;
    END
  END openram_din0[18]
  PIN openram_din0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 296.000 27.050 300.000 ;
    END
  END openram_din0[19]
  PIN openram_din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END openram_din0[1]
  PIN openram_din0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END openram_din0[20]
  PIN openram_din0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 168.680 40.000 169.280 ;
    END
  END openram_din0[21]
  PIN openram_din0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END openram_din0[22]
  PIN openram_din0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 225.800 40.000 226.400 ;
    END
  END openram_din0[23]
  PIN openram_din0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END openram_din0[24]
  PIN openram_din0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 296.000 24.290 300.000 ;
    END
  END openram_din0[25]
  PIN openram_din0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END openram_din0[26]
  PIN openram_din0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END openram_din0[27]
  PIN openram_din0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 273.400 40.000 274.000 ;
    END
  END openram_din0[28]
  PIN openram_din0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 253.000 40.000 253.600 ;
    END
  END openram_din0[29]
  PIN openram_din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 114.280 40.000 114.880 ;
    END
  END openram_din0[2]
  PIN openram_din0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END openram_din0[30]
  PIN openram_din0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END openram_din0[31]
  PIN openram_din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 257.080 40.000 257.680 ;
    END
  END openram_din0[3]
  PIN openram_din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END openram_din0[4]
  PIN openram_din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 145.560 40.000 146.160 ;
    END
  END openram_din0[5]
  PIN openram_din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 248.920 40.000 249.520 ;
    END
  END openram_din0[6]
  PIN openram_din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 175.480 40.000 176.080 ;
    END
  END openram_din0[7]
  PIN openram_din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 296.000 11.410 300.000 ;
    END
  END openram_din0[8]
  PIN openram_din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 296.000 8.650 300.000 ;
    END
  END openram_din0[9]
  PIN openram_dout0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 280.200 40.000 280.800 ;
    END
  END openram_dout0[0]
  PIN openram_dout0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END openram_dout0[10]
  PIN openram_dout0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END openram_dout0[11]
  PIN openram_dout0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 13.640 40.000 14.240 ;
    END
  END openram_dout0[12]
  PIN openram_dout0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 292.440 40.000 293.040 ;
    END
  END openram_dout0[13]
  PIN openram_dout0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END openram_dout0[14]
  PIN openram_dout0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END openram_dout0[15]
  PIN openram_dout0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END openram_dout0[16]
  PIN openram_dout0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 219.000 40.000 219.600 ;
    END
  END openram_dout0[17]
  PIN openram_dout0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 148.280 40.000 148.880 ;
    END
  END openram_dout0[18]
  PIN openram_dout0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END openram_dout0[19]
  PIN openram_dout0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END openram_dout0[1]
  PIN openram_dout0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 55.800 40.000 56.400 ;
    END
  END openram_dout0[20]
  PIN openram_dout0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END openram_dout0[21]
  PIN openram_dout0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 276.120 40.000 276.720 ;
    END
  END openram_dout0[22]
  PIN openram_dout0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 202.680 40.000 203.280 ;
    END
  END openram_dout0[23]
  PIN openram_dout0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END openram_dout0[24]
  PIN openram_dout0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 74.840 40.000 75.440 ;
    END
  END openram_dout0[25]
  PIN openram_dout0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 296.000 14.170 300.000 ;
    END
  END openram_dout0[26]
  PIN openram_dout0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END openram_dout0[27]
  PIN openram_dout0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 296.000 32.570 300.000 ;
    END
  END openram_dout0[28]
  PIN openram_dout0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 125.160 40.000 125.760 ;
    END
  END openram_dout0[29]
  PIN openram_dout0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 296.000 29.810 300.000 ;
    END
  END openram_dout0[2]
  PIN openram_dout0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 156.440 40.000 157.040 ;
    END
  END openram_dout0[30]
  PIN openram_dout0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 24.520 40.000 25.120 ;
    END
  END openram_dout0[31]
  PIN openram_dout0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 195.880 40.000 196.480 ;
    END
  END openram_dout0[3]
  PIN openram_dout0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 296.000 19.690 300.000 ;
    END
  END openram_dout0[4]
  PIN openram_dout0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 78.920 40.000 79.520 ;
    END
  END openram_dout0[5]
  PIN openram_dout0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END openram_dout0[6]
  PIN openram_dout0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END openram_dout0[7]
  PIN openram_dout0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END openram_dout0[8]
  PIN openram_dout0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END openram_dout0[9]
  PIN openram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 210.840 40.000 211.440 ;
    END
  END openram_web0
  PIN openram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END openram_wmask0[0]
  PIN openram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END openram_wmask0[1]
  PIN openram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END openram_wmask0[2]
  PIN openram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 265.240 40.000 265.840 ;
    END
  END openram_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.545 10.640 11.145 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.195 10.640 20.795 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.850 10.640 30.450 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.370 10.640 15.970 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.025 10.640 25.625 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 83.000 40.000 83.600 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 296.000 38.090 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 1.400 40.000 2.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 129.240 40.000 129.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 9.560 40.000 10.160 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 91.160 40.000 91.760 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 51.720 40.000 52.320 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 214.920 40.000 215.520 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 183.640 40.000 184.240 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 296.000 22.450 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 87.080 40.000 87.680 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 288.360 40.000 288.960 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 223.080 40.000 223.680 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 121.080 40.000 121.680 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 229.880 40.000 230.480 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 36.760 40.000 37.360 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 70.760 40.000 71.360 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 110.200 40.000 110.800 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 191.800 40.000 192.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 152.360 40.000 152.960 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 20.440 40.000 21.040 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 269.320 40.000 269.920 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 233.960 40.000 234.560 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 171.400 40.000 172.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 198.600 40.000 199.200 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 133.320 40.000 133.920 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 40.840 40.000 41.440 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 261.160 40.000 261.760 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 179.560 40.000 180.160 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 63.960 40.000 64.560 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 137.400 40.000 138.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 97.960 40.000 98.560 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 16.360 40.000 16.960 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 284.280 40.000 284.880 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 238.040 40.000 238.640 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 106.120 40.000 106.720 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 187.720 40.000 188.320 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 296.000 39.930 300.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 118.360 40.000 118.960 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 296.000 35.330 300.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 47.640 40.000 48.240 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 296.000 1.290 300.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 32.680 40.000 33.280 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 296.000 16.930 300.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 160.520 40.000 161.120 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 246.200 40.000 246.800 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 5.480 40.000 6.080 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 242.120 40.000 242.720 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 43.560 40.000 44.160 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 296.000 5.890 300.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 296.000 4.050 300.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 68.040 40.000 68.640 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 206.760 40.000 207.360 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 4.285 10.795 39.875 296.735 ;
      LAYER met1 ;
        RECT 0.070 10.640 39.950 296.780 ;
      LAYER met2 ;
        RECT 0.100 295.720 0.730 298.365 ;
        RECT 1.570 295.720 3.490 298.365 ;
        RECT 4.330 295.720 5.330 298.365 ;
        RECT 6.170 295.720 8.090 298.365 ;
        RECT 8.930 295.720 10.850 298.365 ;
        RECT 11.690 295.720 13.610 298.365 ;
        RECT 14.450 295.720 16.370 298.365 ;
        RECT 17.210 295.720 19.130 298.365 ;
        RECT 19.970 295.720 21.890 298.365 ;
        RECT 22.730 295.720 23.730 298.365 ;
        RECT 24.570 295.720 26.490 298.365 ;
        RECT 27.330 295.720 29.250 298.365 ;
        RECT 30.090 295.720 32.010 298.365 ;
        RECT 32.850 295.720 34.770 298.365 ;
        RECT 35.610 295.720 37.530 298.365 ;
        RECT 38.370 295.720 39.370 298.365 ;
        RECT 0.100 4.280 39.920 295.720 ;
        RECT 0.650 1.515 1.650 4.280 ;
        RECT 2.490 1.515 4.410 4.280 ;
        RECT 5.250 1.515 7.170 4.280 ;
        RECT 8.010 1.515 9.930 4.280 ;
        RECT 10.770 1.515 12.690 4.280 ;
        RECT 13.530 1.515 15.450 4.280 ;
        RECT 16.290 1.515 17.290 4.280 ;
        RECT 18.130 1.515 20.050 4.280 ;
        RECT 20.890 1.515 22.810 4.280 ;
        RECT 23.650 1.515 25.570 4.280 ;
        RECT 26.410 1.515 28.330 4.280 ;
        RECT 29.170 1.515 31.090 4.280 ;
        RECT 31.930 1.515 33.850 4.280 ;
        RECT 34.690 1.515 35.690 4.280 ;
        RECT 36.530 1.515 38.450 4.280 ;
        RECT 39.290 1.515 39.920 4.280 ;
      LAYER met3 ;
        RECT 4.400 297.520 36.490 298.345 ;
        RECT 4.400 297.480 35.600 297.520 ;
        RECT 3.070 296.120 35.600 297.480 ;
        RECT 3.070 294.800 36.490 296.120 ;
        RECT 4.400 293.440 36.490 294.800 ;
        RECT 4.400 293.400 35.600 293.440 ;
        RECT 3.070 292.040 35.600 293.400 ;
        RECT 3.070 290.720 36.490 292.040 ;
        RECT 4.400 289.360 36.490 290.720 ;
        RECT 4.400 289.320 35.600 289.360 ;
        RECT 3.070 287.960 35.600 289.320 ;
        RECT 3.070 286.640 36.490 287.960 ;
        RECT 4.400 285.280 36.490 286.640 ;
        RECT 4.400 285.240 35.600 285.280 ;
        RECT 3.070 283.920 35.600 285.240 ;
        RECT 4.400 283.880 35.600 283.920 ;
        RECT 4.400 282.520 36.490 283.880 ;
        RECT 3.070 281.200 36.490 282.520 ;
        RECT 3.070 279.840 35.600 281.200 ;
        RECT 4.400 279.800 35.600 279.840 ;
        RECT 4.400 278.440 36.490 279.800 ;
        RECT 3.070 277.120 36.490 278.440 ;
        RECT 3.070 275.760 35.600 277.120 ;
        RECT 4.400 275.720 35.600 275.760 ;
        RECT 4.400 274.400 36.490 275.720 ;
        RECT 4.400 274.360 35.600 274.400 ;
        RECT 3.070 273.000 35.600 274.360 ;
        RECT 3.070 271.680 36.490 273.000 ;
        RECT 4.400 270.320 36.490 271.680 ;
        RECT 4.400 270.280 35.600 270.320 ;
        RECT 3.070 268.920 35.600 270.280 ;
        RECT 3.070 267.600 36.490 268.920 ;
        RECT 4.400 266.240 36.490 267.600 ;
        RECT 4.400 266.200 35.600 266.240 ;
        RECT 3.070 264.840 35.600 266.200 ;
        RECT 3.070 263.520 36.490 264.840 ;
        RECT 4.400 262.160 36.490 263.520 ;
        RECT 4.400 262.120 35.600 262.160 ;
        RECT 3.070 260.760 35.600 262.120 ;
        RECT 3.070 259.440 36.490 260.760 ;
        RECT 4.400 258.080 36.490 259.440 ;
        RECT 4.400 258.040 35.600 258.080 ;
        RECT 3.070 256.720 35.600 258.040 ;
        RECT 4.400 256.680 35.600 256.720 ;
        RECT 4.400 255.320 36.490 256.680 ;
        RECT 3.070 254.000 36.490 255.320 ;
        RECT 3.070 252.640 35.600 254.000 ;
        RECT 4.400 252.600 35.600 252.640 ;
        RECT 4.400 251.240 36.490 252.600 ;
        RECT 3.070 249.920 36.490 251.240 ;
        RECT 3.070 248.560 35.600 249.920 ;
        RECT 4.400 248.520 35.600 248.560 ;
        RECT 4.400 247.200 36.490 248.520 ;
        RECT 4.400 247.160 35.600 247.200 ;
        RECT 3.070 245.800 35.600 247.160 ;
        RECT 3.070 244.480 36.490 245.800 ;
        RECT 4.400 243.120 36.490 244.480 ;
        RECT 4.400 243.080 35.600 243.120 ;
        RECT 3.070 241.720 35.600 243.080 ;
        RECT 3.070 240.400 36.490 241.720 ;
        RECT 4.400 239.040 36.490 240.400 ;
        RECT 4.400 239.000 35.600 239.040 ;
        RECT 3.070 237.640 35.600 239.000 ;
        RECT 3.070 236.320 36.490 237.640 ;
        RECT 4.400 234.960 36.490 236.320 ;
        RECT 4.400 234.920 35.600 234.960 ;
        RECT 3.070 233.560 35.600 234.920 ;
        RECT 3.070 232.240 36.490 233.560 ;
        RECT 4.400 230.880 36.490 232.240 ;
        RECT 4.400 230.840 35.600 230.880 ;
        RECT 3.070 229.520 35.600 230.840 ;
        RECT 4.400 229.480 35.600 229.520 ;
        RECT 4.400 228.120 36.490 229.480 ;
        RECT 3.070 226.800 36.490 228.120 ;
        RECT 3.070 225.440 35.600 226.800 ;
        RECT 4.400 225.400 35.600 225.440 ;
        RECT 4.400 224.080 36.490 225.400 ;
        RECT 4.400 224.040 35.600 224.080 ;
        RECT 3.070 222.680 35.600 224.040 ;
        RECT 3.070 221.360 36.490 222.680 ;
        RECT 4.400 220.000 36.490 221.360 ;
        RECT 4.400 219.960 35.600 220.000 ;
        RECT 3.070 218.600 35.600 219.960 ;
        RECT 3.070 217.280 36.490 218.600 ;
        RECT 4.400 215.920 36.490 217.280 ;
        RECT 4.400 215.880 35.600 215.920 ;
        RECT 3.070 214.520 35.600 215.880 ;
        RECT 3.070 213.200 36.490 214.520 ;
        RECT 4.400 211.840 36.490 213.200 ;
        RECT 4.400 211.800 35.600 211.840 ;
        RECT 3.070 210.440 35.600 211.800 ;
        RECT 3.070 209.120 36.490 210.440 ;
        RECT 4.400 207.760 36.490 209.120 ;
        RECT 4.400 207.720 35.600 207.760 ;
        RECT 3.070 206.400 35.600 207.720 ;
        RECT 4.400 206.360 35.600 206.400 ;
        RECT 4.400 205.000 36.490 206.360 ;
        RECT 3.070 203.680 36.490 205.000 ;
        RECT 3.070 202.320 35.600 203.680 ;
        RECT 4.400 202.280 35.600 202.320 ;
        RECT 4.400 200.920 36.490 202.280 ;
        RECT 3.070 199.600 36.490 200.920 ;
        RECT 3.070 198.240 35.600 199.600 ;
        RECT 4.400 198.200 35.600 198.240 ;
        RECT 4.400 196.880 36.490 198.200 ;
        RECT 4.400 196.840 35.600 196.880 ;
        RECT 3.070 195.480 35.600 196.840 ;
        RECT 3.070 194.160 36.490 195.480 ;
        RECT 4.400 192.800 36.490 194.160 ;
        RECT 4.400 192.760 35.600 192.800 ;
        RECT 3.070 191.400 35.600 192.760 ;
        RECT 3.070 190.080 36.490 191.400 ;
        RECT 4.400 188.720 36.490 190.080 ;
        RECT 4.400 188.680 35.600 188.720 ;
        RECT 3.070 187.320 35.600 188.680 ;
        RECT 3.070 186.000 36.490 187.320 ;
        RECT 4.400 184.640 36.490 186.000 ;
        RECT 4.400 184.600 35.600 184.640 ;
        RECT 3.070 183.240 35.600 184.600 ;
        RECT 3.070 181.920 36.490 183.240 ;
        RECT 4.400 180.560 36.490 181.920 ;
        RECT 4.400 180.520 35.600 180.560 ;
        RECT 3.070 179.200 35.600 180.520 ;
        RECT 4.400 179.160 35.600 179.200 ;
        RECT 4.400 177.800 36.490 179.160 ;
        RECT 3.070 176.480 36.490 177.800 ;
        RECT 3.070 175.120 35.600 176.480 ;
        RECT 4.400 175.080 35.600 175.120 ;
        RECT 4.400 173.720 36.490 175.080 ;
        RECT 3.070 172.400 36.490 173.720 ;
        RECT 3.070 171.040 35.600 172.400 ;
        RECT 4.400 171.000 35.600 171.040 ;
        RECT 4.400 169.680 36.490 171.000 ;
        RECT 4.400 169.640 35.600 169.680 ;
        RECT 3.070 168.280 35.600 169.640 ;
        RECT 3.070 166.960 36.490 168.280 ;
        RECT 4.400 165.600 36.490 166.960 ;
        RECT 4.400 165.560 35.600 165.600 ;
        RECT 3.070 164.200 35.600 165.560 ;
        RECT 3.070 162.880 36.490 164.200 ;
        RECT 4.400 161.520 36.490 162.880 ;
        RECT 4.400 161.480 35.600 161.520 ;
        RECT 3.070 160.120 35.600 161.480 ;
        RECT 3.070 158.800 36.490 160.120 ;
        RECT 4.400 157.440 36.490 158.800 ;
        RECT 4.400 157.400 35.600 157.440 ;
        RECT 3.070 156.040 35.600 157.400 ;
        RECT 3.070 154.720 36.490 156.040 ;
        RECT 4.400 153.360 36.490 154.720 ;
        RECT 4.400 153.320 35.600 153.360 ;
        RECT 3.070 152.000 35.600 153.320 ;
        RECT 4.400 151.960 35.600 152.000 ;
        RECT 4.400 150.600 36.490 151.960 ;
        RECT 3.070 149.280 36.490 150.600 ;
        RECT 3.070 147.920 35.600 149.280 ;
        RECT 4.400 147.880 35.600 147.920 ;
        RECT 4.400 146.560 36.490 147.880 ;
        RECT 4.400 146.520 35.600 146.560 ;
        RECT 3.070 145.160 35.600 146.520 ;
        RECT 3.070 143.840 36.490 145.160 ;
        RECT 4.400 142.480 36.490 143.840 ;
        RECT 4.400 142.440 35.600 142.480 ;
        RECT 3.070 141.080 35.600 142.440 ;
        RECT 3.070 139.760 36.490 141.080 ;
        RECT 4.400 138.400 36.490 139.760 ;
        RECT 4.400 138.360 35.600 138.400 ;
        RECT 3.070 137.000 35.600 138.360 ;
        RECT 3.070 135.680 36.490 137.000 ;
        RECT 4.400 134.320 36.490 135.680 ;
        RECT 4.400 134.280 35.600 134.320 ;
        RECT 3.070 132.920 35.600 134.280 ;
        RECT 3.070 131.600 36.490 132.920 ;
        RECT 4.400 130.240 36.490 131.600 ;
        RECT 4.400 130.200 35.600 130.240 ;
        RECT 3.070 128.880 35.600 130.200 ;
        RECT 4.400 128.840 35.600 128.880 ;
        RECT 4.400 127.480 36.490 128.840 ;
        RECT 3.070 126.160 36.490 127.480 ;
        RECT 3.070 124.800 35.600 126.160 ;
        RECT 4.400 124.760 35.600 124.800 ;
        RECT 4.400 123.400 36.490 124.760 ;
        RECT 3.070 122.080 36.490 123.400 ;
        RECT 3.070 120.720 35.600 122.080 ;
        RECT 4.400 120.680 35.600 120.720 ;
        RECT 4.400 119.360 36.490 120.680 ;
        RECT 4.400 119.320 35.600 119.360 ;
        RECT 3.070 117.960 35.600 119.320 ;
        RECT 3.070 116.640 36.490 117.960 ;
        RECT 4.400 115.280 36.490 116.640 ;
        RECT 4.400 115.240 35.600 115.280 ;
        RECT 3.070 113.880 35.600 115.240 ;
        RECT 3.070 112.560 36.490 113.880 ;
        RECT 4.400 111.200 36.490 112.560 ;
        RECT 4.400 111.160 35.600 111.200 ;
        RECT 3.070 109.800 35.600 111.160 ;
        RECT 3.070 108.480 36.490 109.800 ;
        RECT 4.400 107.120 36.490 108.480 ;
        RECT 4.400 107.080 35.600 107.120 ;
        RECT 3.070 105.720 35.600 107.080 ;
        RECT 3.070 104.400 36.490 105.720 ;
        RECT 4.400 103.040 36.490 104.400 ;
        RECT 4.400 103.000 35.600 103.040 ;
        RECT 3.070 101.680 35.600 103.000 ;
        RECT 4.400 101.640 35.600 101.680 ;
        RECT 4.400 100.280 36.490 101.640 ;
        RECT 3.070 98.960 36.490 100.280 ;
        RECT 3.070 97.600 35.600 98.960 ;
        RECT 4.400 97.560 35.600 97.600 ;
        RECT 4.400 96.200 36.490 97.560 ;
        RECT 3.070 94.880 36.490 96.200 ;
        RECT 3.070 93.520 35.600 94.880 ;
        RECT 4.400 93.480 35.600 93.520 ;
        RECT 4.400 92.160 36.490 93.480 ;
        RECT 4.400 92.120 35.600 92.160 ;
        RECT 3.070 90.760 35.600 92.120 ;
        RECT 3.070 89.440 36.490 90.760 ;
        RECT 4.400 88.080 36.490 89.440 ;
        RECT 4.400 88.040 35.600 88.080 ;
        RECT 3.070 86.680 35.600 88.040 ;
        RECT 3.070 85.360 36.490 86.680 ;
        RECT 4.400 84.000 36.490 85.360 ;
        RECT 4.400 83.960 35.600 84.000 ;
        RECT 3.070 82.600 35.600 83.960 ;
        RECT 3.070 81.280 36.490 82.600 ;
        RECT 4.400 79.920 36.490 81.280 ;
        RECT 4.400 79.880 35.600 79.920 ;
        RECT 3.070 78.520 35.600 79.880 ;
        RECT 3.070 77.200 36.490 78.520 ;
        RECT 4.400 75.840 36.490 77.200 ;
        RECT 4.400 75.800 35.600 75.840 ;
        RECT 3.070 74.480 35.600 75.800 ;
        RECT 4.400 74.440 35.600 74.480 ;
        RECT 4.400 73.080 36.490 74.440 ;
        RECT 3.070 71.760 36.490 73.080 ;
        RECT 3.070 70.400 35.600 71.760 ;
        RECT 4.400 70.360 35.600 70.400 ;
        RECT 4.400 69.040 36.490 70.360 ;
        RECT 4.400 69.000 35.600 69.040 ;
        RECT 3.070 67.640 35.600 69.000 ;
        RECT 3.070 66.320 36.490 67.640 ;
        RECT 4.400 64.960 36.490 66.320 ;
        RECT 4.400 64.920 35.600 64.960 ;
        RECT 3.070 63.560 35.600 64.920 ;
        RECT 3.070 62.240 36.490 63.560 ;
        RECT 4.400 60.880 36.490 62.240 ;
        RECT 4.400 60.840 35.600 60.880 ;
        RECT 3.070 59.480 35.600 60.840 ;
        RECT 3.070 58.160 36.490 59.480 ;
        RECT 4.400 56.800 36.490 58.160 ;
        RECT 4.400 56.760 35.600 56.800 ;
        RECT 3.070 55.400 35.600 56.760 ;
        RECT 3.070 54.080 36.490 55.400 ;
        RECT 4.400 52.720 36.490 54.080 ;
        RECT 4.400 52.680 35.600 52.720 ;
        RECT 3.070 51.360 35.600 52.680 ;
        RECT 4.400 51.320 35.600 51.360 ;
        RECT 4.400 49.960 36.490 51.320 ;
        RECT 3.070 48.640 36.490 49.960 ;
        RECT 3.070 47.280 35.600 48.640 ;
        RECT 4.400 47.240 35.600 47.280 ;
        RECT 4.400 45.880 36.490 47.240 ;
        RECT 3.070 44.560 36.490 45.880 ;
        RECT 3.070 43.200 35.600 44.560 ;
        RECT 4.400 43.160 35.600 43.200 ;
        RECT 4.400 41.840 36.490 43.160 ;
        RECT 4.400 41.800 35.600 41.840 ;
        RECT 3.070 40.440 35.600 41.800 ;
        RECT 3.070 39.120 36.490 40.440 ;
        RECT 4.400 37.760 36.490 39.120 ;
        RECT 4.400 37.720 35.600 37.760 ;
        RECT 3.070 36.360 35.600 37.720 ;
        RECT 3.070 35.040 36.490 36.360 ;
        RECT 4.400 33.680 36.490 35.040 ;
        RECT 4.400 33.640 35.600 33.680 ;
        RECT 3.070 32.280 35.600 33.640 ;
        RECT 3.070 30.960 36.490 32.280 ;
        RECT 4.400 29.600 36.490 30.960 ;
        RECT 4.400 29.560 35.600 29.600 ;
        RECT 3.070 28.200 35.600 29.560 ;
        RECT 3.070 26.880 36.490 28.200 ;
        RECT 4.400 25.520 36.490 26.880 ;
        RECT 4.400 25.480 35.600 25.520 ;
        RECT 3.070 24.160 35.600 25.480 ;
        RECT 4.400 24.120 35.600 24.160 ;
        RECT 4.400 22.760 36.490 24.120 ;
        RECT 3.070 21.440 36.490 22.760 ;
        RECT 3.070 20.080 35.600 21.440 ;
        RECT 4.400 20.040 35.600 20.080 ;
        RECT 4.400 18.680 36.490 20.040 ;
        RECT 3.070 17.360 36.490 18.680 ;
        RECT 3.070 16.000 35.600 17.360 ;
        RECT 4.400 15.960 35.600 16.000 ;
        RECT 4.400 14.640 36.490 15.960 ;
        RECT 4.400 14.600 35.600 14.640 ;
        RECT 3.070 13.240 35.600 14.600 ;
        RECT 3.070 11.920 36.490 13.240 ;
        RECT 4.400 10.560 36.490 11.920 ;
        RECT 4.400 10.520 35.600 10.560 ;
        RECT 3.070 9.160 35.600 10.520 ;
        RECT 3.070 7.840 36.490 9.160 ;
        RECT 4.400 6.480 36.490 7.840 ;
        RECT 4.400 6.440 35.600 6.480 ;
        RECT 3.070 5.080 35.600 6.440 ;
        RECT 3.070 3.760 36.490 5.080 ;
        RECT 4.400 2.400 36.490 3.760 ;
        RECT 4.400 2.360 35.600 2.400 ;
        RECT 3.070 1.535 35.600 2.360 ;
      LAYER met4 ;
        RECT 5.815 10.240 9.145 288.560 ;
        RECT 11.545 10.240 13.970 288.560 ;
        RECT 16.370 10.240 18.795 288.560 ;
        RECT 5.815 6.975 20.800 10.240 ;
  END
END wrapped_wb_openram_shim
END LIBRARY

